module vnds

pub enum BgType as u32
{
	text8bpp
	text4bpp
	rotation
	exrotation
	bmp8
	bmp16
}

pub enum BgSize as u32
{
	r_128x128 =   (0 << 14) 
	r_256x256 =   (1 << 14) 
	r_512x512 =   (2 << 14) 
	r_1024x1024 = (3 << 14) 
	
	t_256x256 = (0 << 14) | (1 << 16)
	t_512x256 = (1 << 14) | (1 << 16)
	t_256x512 = (2 << 14) | (1 << 16)
	t_512x512 = (3 << 14) | (1 << 16)
	
	er_128x128 = (0 << 14) | (2 << 16)
	er_256x256 = (1 << 14) | (2 << 16)
	er_512x512 = (2 << 14) | (2 << 16)
	er_1024x1024 = (3 << 14) | (2 << 16)
	
	b8_128x128 =  ((0 << 14) | (1 << 7) | (3 << 16))
	b8_256x256 =  ((1 << 14) | (1 << 7) | (3 << 16))
	b8_512x256 =  ((2 << 14) | (1 << 7) | (3 << 16))
	b8_512x512 =  ((3 << 14) | (1 << 7) | (3 << 16))
	b8_1024x512 = ((1 << 14) | (3 << 16))
	b8_512x1024 = ((0      ) | (3 << 16))
	b16_128x128 = ((0 << 14) | (1 << 7) | (1 << 2) | (4 << 16))
	b16_256x256 = ((1 << 14) | (1 << 7) | (1 << 2) | (4 << 16))
	b16_512x256 = ((2 << 14) | (1 << 7) | (1 << 2) | (4 << 16))
	b16_512x512 = ((3 << 14) | (1 << 7) | (1 << 2) | (4 << 16))
}